/home/linux/ieng6/ee260bwi20/kexia/lab3/libdir/lef/tcbn65gplus_8lmT2.lef